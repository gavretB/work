module imem(cur_addr, inst);
input [11:0] cur_addr;
output [18:0] inst;

function [18:0] dec;
input [11:0] in;
	case(in)
/*
	//test.ppe
		0: dec = 19'b1110000000000010000;	// jmp	16
		1: dec = 19'b1001011100000000000; // inp	r7, 0(r0)
		2: dec = 19'b1000011000000000000;	// ldm	r6, 0(r0)
		3: dec = 19'b1000111111000000001; // stm	r7, 1(r6)
		4: dec = 19'b0100111011000000001; // add	r6, r6, 1
		5: dec = 19'b1000111000000000000; // stm	r6, 0(r0)
		6: dec = 19'b1111010000000000000; // reti
		16: dec = 19'b1111100000000000000; // enai -> 割り込み受付る
		17: dec = 19'b1000001100000000000; // ldm	r3, 0(r0) -> r3:dmem(r0+0)
		18: dec = 19'b0001001101101000000; // sub	r3, r3, r2 -> r3: r3-r2
		19: dec = 19'b1010000000011111101; // bz	-3 -> 17へ
		20: dec = 19'b1000001101000000001; // ldm	r3, 1(r2) -> r3: dmem(r2+1)
		21: dec = 19'b1001101100000001111; // out	r3, 15(r0)
		22: dec = 19'b0100001001000000001; // add	r2, r2, 1 -> r2 = r2 + 1
		23: dec = 19'b1110000000000010001; // jmp	17
		default:dec=19'b0000000000000000000;
*/
/*
		0:16行目へ
		16:割り込みを受け入れ設定
		17:r3にdmem（r0+0）を書き出し
		18:r3にr3-r2を代入
		19:17行目へ
		....
		割り込み発生で1へ
		1:r7をdmem(r0+0)へ
		2:dmem(r0+0)をr6へ
		3:r7をdmem(r6+1)へ
		4:r6+1=r6へ
		5:r6をdmem(r0+0)へ
		6:割り込み発生アドレスの次のアドレスへ
*/

/*	//test1A.ppe
		0: dec = 19'b1110000000000010000;	// jmp	16
		1: dec = 19'b1111010000000000000; // reti
		16: dec = 19'b1111100000000000000;	// enai
		17: dec = 19'b0100000100000001010; // add r1, r0, 10
		18: dec = 19'b1000100100000000000; // stm	r1, 0(r0)
		19: dec = 19'b0101000100100000001; // sub	r1, r1, 1
		20: dec = 19'b1010100000011111101; //	bnz	-3
		21: dec = 19'b1110000000000010101; //	jmp	21
*/
/*
		0:16行目へ
		16:割り込みを受け入れ設定
		17:r1 = r0 + 10 = 0 + 10 = 10
		18:dmem(r0+0) = r1 -> dmem[0] = 10
		19:r1 = r1-1 = 10 - 1 = 9
		20:18へ
		18:dmem(r0+0) = r1 -> dmem[0] = 9
		19:r1 = 8
		20:18へ
		...
		r1=0のとき
		20:21へ
		21:18へ
		18:dmem[0] = 0
		...
		20:
*/
/*
 //mem_IO挙動確認コード
		0: dec = 19'b0100000100000001010; // add	r1, r0, 10
		1: dec = 19'b0100001000000010000; // add	r2, r0, 16
		2: dec = 19'b1000100101000000000; //	stm	r1, 0(r2)
		3: dec = 19'b1000000101000000001; // ldm	r1, 1(r2)
		4: dec = 19'b1110000000000000000; //	jmp	0
*/
/*
	//test1B.ppe
		0: dec = 19'b1110000000000010000; //	jmp	16
		1: dec = 19'b1000011101000000000; //	ldm	r7, 0(r2)
		2: dec = 19'b0101011111100000001; //	sub	r7, r7, 1
		3: dec = 19'b1000111101000000000; //	stm	r7, 0(r2)
		4: dec = 19'b1111010000000000000; //	reti
		16: dec = 19'b1111110000000000000; //	disi
		17: dec = 19'b0100001000000010000; // add	r2, r0, 16
		18: dec = 19'b0100000100000001010; // add	r1, r0, 10
		19: dec = 19'b1000100101000000000; //	stm	r1, 0(r2)
		20: dec = 19'b1111100000000000000; //	enai
		21: dec = 19'b1000000101000000000; // ldm	r1, 0(r2)
		22: dec = 19'b0100000100100000000; //	add	r1, r1, r0
		23: dec = 19'b1010100000011111101; //	bnz	-3
		24: dec = 19'b1110000000000011000; //	jmp	24
*/
/*
		0:16行目へ
		16:割り込みを拒否設定
		17:r2 = r0 + 16 = 16
		18:r1 = r0 + 10 = 10
		19:dmem(r2+0) = r1 = dmem[16] = 10
		20:割り込みを受諾設定
		21:r1 = dmem[r2+0] = dmem[16] = 10
		22:r1 = r1 + r0 = 10
		23:21へ
		21:r1 = dmem[r2+0] = dmem[16] = 10
		...
		割り込み
		1:r7 = dmem[r2+0] = dmem[16] = 10
		2:r7 = 9
		3:dmem[16] = 9
*/
/*
//test2.ppe
	0: dec = 19'b1110000000000010000; //	jmp	16
	1: dec = 19'b1111010000000000000; //	reti
	16: dec = 19'b1111110000000000000; //	disi
	17: dec = 19'b0100100100001111111; //	addc r1, r0, 127
	18: dec = 19'b0100101000110000000; //	addc r2, r1, 128
	19: dec = 19'b0100101101000000001; //	addc r3, r2, 1
	20: dec = 19'b0101110001100000001; //	subc r4, r3, 1
	21: dec = 19'b0101110110010000000; //	subc r5, r4, 128
	22: dec = 19'b0101111010101111101; //	subc r6, r5, 125
	23: dec = 19'b1110000000000010111; //	jmp 23
*/
/*
	0: 16へ
	16: 割り込み拒否
	17: r1 = r0 + 127 = 127, cc_c:0, cc_z:0
	18: r2 = r1 + 128 = 127 + (-128) = -1, cc_c:0, cc_z:0
	19: r3 = r2 + 1 = -1 + 1 = 0, cc_c:0, cc_z:1
	20: r4 = r3 - 1 = 0 - 1 = -1, cc_c:0, cc_z:0
	21: r5 = r4 - (-128) = -1 - (-128) = 127, cc_c:0, cc_z:0
	22: r6 = r5 - 125 = 127 - 125 = 2, cc_c:0, cc_z:0
	23: 23へ
*/
/*
0:dec=19'b1110000000000010000; //	jmp	16
1:dec=19'b1111010000000000000; //	reti
16:dec=19'b1111110000000000000; //	disi
17:dec=19'b0100000100000000001; //	add r1, r0, 1
18:dec=19'b0100001000000000100; //	add r2, r0, 4
19:dec=19'b0100001100000010000; //	add r3, r0, 16
20:dec=19'b0100010000001000000; //	add r4, r0, 64
21:dec=19'b0001010101110000000; //	sub r5, r3, r4
default:dec=19'b0000000000000000000;
*/
/*
//test3.ppe
	0:dec=19'b1110000000000010000; //	jmp	16
	1:dec=19'b1111010000000000000; //	reti
	16:dec=19'b1111110000000000000; //	disi
	17:dec=19'b0100000100000000001; //	add r1, r0, 1
	18:dec=19'b0100001000000000100; //	add r2, r0, 4
	19:dec=19'b0100001100000010000; //	add r3, r0, 16
	20:dec=19'b0100010000001000000; //	add r4, r0, 64
	21:dec=19'b0000010100000000000; //	add r5, r0, r0
	22:dec=19'b0010110110100100000; // 	or  r5, r5, r1
	23:dec=19'b0010110110101000000; // 	or  r5, r5, r2
	24:dec=19'b0010110110101100000; // 	or  r5, r5, r3
	25:dec=19'b0010110110110000000; // 	or  r5, r5, r4

	26:dec=19'b1100000100100100000; // 	shl r1, r1, 1
	27:dec=19'b1100001001000100000; // 	shl r2, r2, 1
	28:dec=19'b1100001101100100000; // 	shl r3, r3, 1
	29:dec=19'b1100010010000100000; //	shl r4, r4, 1
	30:dec=19'b0010110110100100000; //	or  r5, r5, r1
	31:dec=19'b0010110110101000000; //	or  r5, r5, r2
	32:dec=19'b0010110110101100000; //	or  r5, r5, r3
	33:dec=19'b0010110110110000000; //	or  r5, r5, r4

	34:dec=19'b1101100100100100011; //	ror r1, r1, 3
	35:dec=19'b1101101001000100011; //	ror r2, r2, 3
	36:dec=19'b1101101101100100011; //	ror r3, r3, 3
	37:dec=19'b1101110010000100011; //	ror r4, r4, 3
	38:dec=19'b0011011010100100000; //	xor r6, r5, r1
	39:dec=19'b0011011011001000000; // 	xor r6, r6, r2
	40:dec=19'b0011011011001100000; // 	xor r6, r6, r3
	41:dec=19'b0011011011010000000; // 	xor r6, r6, r4

	42:dec=19'b0011111110111000000; //	msk r7, r5, r6
	43:dec=19'b0011011111100100000; //	xor r7, r7, r1
	44:dec=19'b0011011111101000000; // 	xor r7, r7, r2
	45:dec=19'b0011011111101100000; // 	xor r7, r7, r3
	46:dec=19'b0011011111110000000; // 	xor r7, r7, r4

	47:dec=19'b1110000000000101111; //	jmp 47
	default:dec=19'b0000000000000000000;
*/
/*
	0: 16へ
	16: 割り込み拒否
	17: r1 = r0 + 1 = 1
	18: r2 = r0 + 4 = 4
	19: r3 = r0 + 16 = 16
	20: r4 = r0 + 64 = 64
	21: r5 = r0 + r0 = 0
	22: r5 = r5 or r1 = 0 or 1 = 1
	23: r5 = r5 or r2 = 1 or 4 = 5
	24: r5 = r5 or r3 = 5 or 16 = 21
	25: r5 = r5 or r4 = 21 or 64 = 00010101 or 01000000 = 01010101 = 85
	26: r1 = r1 shl 1 = 1 shl 1 = 2
	27: r2 = r2 shl 1 = 4 shl 1 = 8
	28: r3 = r3 shl 1 = 16 shl 1 = 32
	29: r4 = r4 shl 1 = 64 shl 1 = 128
	30: r5 = r5 or r1 = 85 or 2 = 01010101 or 00000010 = 01010111 = 87
	31: r5 = r5 or r2 = 87 or 8 = 01010111 or 00001000 = 01011111 = 95
	32: r5 = r5 or r3 = 95 or 32 = 01011111 or 00100000 = 01111111 = 127
	33: r5 = r5 or r4 = 127 or 128 = 255
	34: r1 =r1 ror 3 = 2 ror 3 = 00000010 ror 3 = 01000000 = 64
	35: r2 = r2 ror 3 = 8 ror 3 = 00001000 ror 3 = 00000001 = 1
	36: r3 = r3 ror 3 = 32 ror 3 = 00100000 ror 3 = 00000100 = 4
	37: r4 = r4 ror 3 = 128 ror 3 = 10000000 ror 3 = 00010000 = 16
	38: r6 = r5 xor r1 = 255 xor 64 = 11111111 xor 01000000 = 10111111 = 255-64=191
	39: r6 = r6 xor r2 = 191 xor 1 = 10111111 xor 00000001 = 10111110 = 190
	40: r6 = r6 xor r3 = 190 xor 4 = 10111110 xor 00000100 = 10111010 = 186
	41: r6 = r6 xor r4 = 186 xor 16 = 10111010 xor 00010000 = 10101010 = 170
	42: r7 = r5 msk r6 = 255 msk 170 = 11111111 msk 10101010 = 01010101 = 64 + 16 + 4 + 1 = 85
	43: r7 = r7 xor r1 = 85 xor 64 = 01010101 xor 01000000 = 00010101 = 21
	44: r7 = r7 xor r2 = 21 xor 1 = 00010101 xor 00000001 = 00010100 = 20
	45: r7 = r7 xor r3 = 20 xor 4 = 00010100 xor 00000100 = 00010000 = 16
	46: r7 = r7 xor r4 = 16 xor 16 = 00010000 xor 00010000 = 00000000 = 0
	47: 47へ
*/
/*
//test4A.ppe
	0:dec=19'b1110000000000010000; //	jmp	16

	1:dec=19'b1111010000000000000; //	reti

	16:dec=19'b1111100000000000000; //	enai
	17:dec=19'b1001100100000001111; //	out	r1, 15(r0)
	18:dec=19'b0100000100100000001; //	add	r1, r1, 1
	19:dec=19'b0101000000100001010; //	sub	r0, r1, 10
	20:dec=19'b1010100000011111100; //	bnz	-4
	21:dec=19'b1110000000000010101; //	jmp	21
*/
/*
	0:16へ
	16:割り込み受け入れ設定
	17:なし
	18:r1 = r1 + 1 = 0 + 1 = 1
	19:r0 = r1 - 10 = -9
	20:17へ
	21:21へ
*/
/*
//test4B.ppe
	0:dec=19'b1110000000000010000; //	jmp	16

	1:dec=19'b1001011100000000000; //	inp	r7, 0(r0)
	2:dec=19'b1000011000000000000; //	ldm	r6, 0(r0)
	3:dec=19'b1000111111000000001; //	stm	r7, 1(r6)
	4:dec=19'b0100111011000000001; //	add	r6, r6, 1
	5:dec=19'b1000111000000000000; //	stm	r6, 0(r0)
	6:dec=19'b1111010000000000000; //	reti

	16:dec=19'b1111100000000000000; //	enai

	17:dec=19'b1000001100000000000; //	ldm	r3, 0(r0)
	18:dec=19'b0001001101101000000; //	sub	r3, r3, r2
	19:dec=19'b1010000000011111101; //	bz	-3

	20:dec=19'b1000001101000000001; //	ldm	r3, 1(r2)
	21:dec=19'b1001101100000001111; //  out	r3, 15(r0)
	22:dec=19'b0100001001000000001; //	add	r2, r2, 1
	23:dec=19'b1110000000000010001; //	jmp	17
*/
/*
	0:16へ
	16:割り込み受け入れ設定
	17:r3 = dmem(r0+0) = dmem(0) = x
	18:r3 = x - r2 = x - 0 = x
	19:17へ
	20:r3 = dmem(r2+1) = dmem(0+1) = x
	21:なし
	22:r2 = r2 + 1 = 0 + 1 = 1
	23:17へ

	割り込み時
	1:なし
	2:r6 = dmem(r0+0)
	3:dmem(r6+1) = r7
	4:r6 = r6 + 1
	5:dmem(r0+0) = r6
	6:もとアドレスへ
*/

//test5.ppe
	0:dec=19'b1110000000000010000; //	jmp	16

	1:dec=19'b1111010000000000000; //	reti
	2:dec=19'b1000111000011111111; //	stm	r6, 255(r0)
	3:dec=19'b0000011000000000000; //	add	r6, r0, r0
	4:dec=19'b0000011000000000000; //	add	r6, r0, r0
	5:dec=19'b0000000010100000000; //	add	r0, r5, r0
	6:dec=19'b1010000000000000100; //	bz	4

	7:dec=19'b0000011111110000000; //	add	r7, r7, r4
	8:dec=19'b0100111011000000000; //	addc	r6, r6, 0
	9:dec=19'b0101010110100000001; //	sub	r5, r5, 1
	10:dec=19'b1010100000011111100; //	bnz	-4

	11:dec=19'b1000010100011111111; //	ldm	r5, 255(r0)
	12:dec=19'b1000111010100000000; //	stm	r6, 0(r5)
	13:dec=19'b1000111110100000001; //	stm	r7, 1(r5)
	14:dec=19'b1111000000000000000; //	ret

	16:dec=19'b1111110000000000000; //	disi
	17:dec=19'b0100000100000001111; //	add	r1, r0, 15
	18:dec=19'b0100001000000000100; //	add	r2, r0, 4
	19:dec=19'b0100001100000000001; //	add	r3, r0, 1
	20:dec=19'b1000101100000000001; //	stm	r3, 1(r0)
	21:dec=19'b0100001100000000010; //	add	r3, r0, 2
	22:dec=19'b1000101100000000011; //	stm	r3, 3(r0)
	23:dec=19'b0100010000000000011; //	add	r4, r0, 3

	24:dec=19'b0000010101100000000; //	add	r5, r3, r0
	25:dec=19'b0000011001000000000; //	add	r6, r2, r0
	26:dec=19'b1110100000000000010; //	jsb	2
	27:dec=19'b0000001110000000000; //	add	r3, r4, r0
	28:dec=19'b0100010010000000001; //	add	r4, r4, 1
	29:dec=19'b0100001001000000010; //	add	r2, r2, 2
	30:dec=19'b0101000100100000001; //	sub	r1, r1, 1
	31:dec=19'b1010100000011111000; //	bnz	-8

	32:dec=19'b1110000000000100000; //	jmp	32
	default:dec=19'b0000000000000000000;

/*
	0:16へ
	1:reti

	16:disi
	17:add	r1, r0, 15 -> r1 = r0 + 15 = 15
	18:add	r2, r0, 4 -> r2 = r0 + 4 = 4
	19:add	r3, r0, 1 -> r3 = r0 + 1 = 1
	20:stm	r3, 1(r0) -> dmem(r0+1) = r3 = 1
	21:add	r3, r0, 2 -> r3 = r0 + 2 = 2
	22:stm	r3, 3(r0) -> dmem(r0+3) = r3 = 2
	23:add	r4, r0, 3 -> r4 = r0 + 3 = 3

	24:add	r5, r3, r0 -> r5 = r3 + r0 = 2
	25:add	r6, r2, r0 -> r6 = r2 + r0 = 4
	26:jsb	2

	2:stm	r6, 255(r0) -> dmem(r0+255) = r6 = 4
	3:add	r6, r0, r0 -> r6 = r0 + r0 = 0
	4:add	r6, r0, r0 -> r6 = r0 + r0 = 0
	5:add	r0, r5, r0 -> r0 = r5 + r0 = 0
	6:bz	4 -> 11へ

	11:ldm	r5, 255(r0) -> r5 = dmem(r0+255) = x
	12:stm	r6, 0(r5) -> dmem(r5+0) = r6 = 0
	13:stm	r7, 1(r5) -> dmem(r5+1) = r7 =0
	14:ret

	27:add	r3, r4, r0 -> r3 = r4 + r0 =3
	28:add	r4, r4, 1 = r4 = r4 + 1 = 4
	29:add	r2, r2, 2 = 6
	30:sub	r1, r1, 1 = r1 = r1 - 1 = 15 - 1 = 14
	31:bnz	-8 - > 24へ

	32:jmp	32
*/

	endcase
endfunction

assign inst = dec(cur_addr);

endmodule
